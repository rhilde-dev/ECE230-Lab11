module t_flipflop(
    input t,
    input store,
    output memory,
    output n_mem
);

    wire data;
    wire Q, notQ;
    
    multiplexer mux (.A(Q),.B(notQ),.Enable(1'b1), .Sel(t), .Y(data));
    
//    assign data = (j & notQ)|(~k & Q);
    
    d_flipflop dflip (.data(data), .store(store), .memory(Q), .n_mem(notQ));
    
    assign memory = Q;
    assign n_mem = notQ;

endmodule