module jk_flipflop(
    input j,k,
    input store,
    output memory,
    output n_mem
);

    wire data;
    wire Q, notQ;
    
    assign data = (j & notQ)|(~k & Q);
    
    d_flipflop dflip (.data(data), .store(store), .memory(Q), .n_mem(notQ));
    
    assign memory = Q;
    assign n_mem = notQ;

endmodule